module switch_mcu_spi2ahb (
    in_clk  ,
    in_rst  ,
    in_spi_clk,

    
);
// Global signals
input  wire in_clk                   ;
input  wire in_rst                   ;
input  wire in_spi_clk               ;
    
endmodule